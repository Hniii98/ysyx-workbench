`ifndef _MUXKEY_V_
`define _MUXKEY_V_ 

module MuxKey #(
  parameter NR_KEY = 2, 
  parameter KEY_LEN = 1,
  parameter DATA_LEN = 1
) (
  output [DATA_LEN-1:0] out,
  input [KEY_LEN-1:0] key,
  input [NR_KEY*(KEY_LEN + DATA_LEN)-1:0] lut
);
  MuxKeyInternal #(NR_KEY, KEY_LEN, DATA_LEN, 0) i0 (out, key, {DATA_LEN{1'b0}}, lut); // set default to all zero
endmodule

`endif
